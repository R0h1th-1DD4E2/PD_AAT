module round(
)
  
